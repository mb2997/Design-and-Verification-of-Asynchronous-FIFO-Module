// `define WCLK_FRQ 80						//Unit: MHz
// `define RCLK_FRQ 50						//Unit: MHz
// `define WCLK_T/2 ((1/`WCLK_FRQ)/2)
// `define RCLK_T/2 ((1/`RCLK_FRQ)/2)
// `define ADDR_WIDTH 8
// `define DATA_WIDTH 32